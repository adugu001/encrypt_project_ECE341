-- empty for now, but we need a main controller